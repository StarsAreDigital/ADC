module Control (
	input [5:0] ctrl_i,
	output reg memToReg_o,
	output reg memToRead_o,
	output reg memToWrite_o,
	output reg [1:0] aluOp_o,
	output reg regWrite_o
);
	always @(*) begin
		case (ctrl_i)
			6'b000000: begin // Tipo R
				memToReg_o = 1'b0;
				memToRead_o = 1'b0;
				memToWrite_o = 1'b0;
				aluOp_o = 2'b10;
				regWrite_o = 1'b1;
			end
			default: begin
				
			end
		endcase
	end
endmodule
