module REGBANK (
	input [16:0] in,
	output [31:0] out
);
	

endmodule
