module MemWBuffer ( // Memory Access/Write Back
    
);
    
endmodule